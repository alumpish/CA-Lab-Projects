module Ins_Mem (
    input [31:0] in,
    output [31:0] out
  );

  reg [31:0] mem[6:0];

  initial
  begin
    mem[0] = 32'b000000_00001_00010_00000_00000000000;
    mem[1] = 32'b000000_00011_00100_00000_00000000000;
    mem[2] = 32'b000000_00101_00110_00000_00000000000;
    mem[3] = 32'b000000_00111_01000_00010_00000000000;
    mem[4] = 32'b000000_01001_01010_00011_00000000000;
    mem[5] = 32'b000000_01011_01100_00000_00000000000;
    mem[6] = 32'b000000_01101_01110_00000_00000000000;
  end

  assign out = mem[in>>2];

endmodule
